module lexer

[export: 'do_cool_stuff']
fn do_cool_stuff() {
    println('hello from v!')
}

